library verilog;
use verilog.vl_types.all;
entity leitor_txt_vlg_vec_tst is
end leitor_txt_vlg_vec_tst;
