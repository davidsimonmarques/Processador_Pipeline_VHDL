library verilog;
use verilog.vl_types.all;
entity mult4_vlg_vec_tst is
end mult4_vlg_vec_tst;
