library verilog;
use verilog.vl_types.all;
entity ALU_decoder_vlg_vec_tst is
end ALU_decoder_vlg_vec_tst;
