library verilog;
use verilog.vl_types.all;
entity banco_reg_vlg_vec_tst is
end banco_reg_vlg_vec_tst;
