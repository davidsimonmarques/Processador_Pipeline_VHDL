library verilog;
use verilog.vl_types.all;
entity Data_mem_vlg_vec_tst is
end Data_mem_vlg_vec_tst;
