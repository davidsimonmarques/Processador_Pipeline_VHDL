library ieee;
use ieee.std_logic_1164.all;

entity Processador_Pipeline is 

end Processador_Pipeline;

architecture arch_Processador of Processador_Pipeline is
begin

end arch_Processador;