library verilog;
use verilog.vl_types.all;
entity leitor_txt_vlg_check_tst is
    port(
        dataout         : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end leitor_txt_vlg_check_tst;
