library verilog;
use verilog.vl_types.all;
entity Mem_Instr_vlg_vec_tst is
end Mem_Instr_vlg_vec_tst;
